`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
//////////////////////////////////////////////////////////////////////////////////

           
module SE#(WL = 32, INW = 16)
        (input signed [INW-1:0] Imm,
         output signed [WL-1:0] SImm);

assign SImm = { {(WL-INW){Imm[INW-1]}} ,Imm[INW-1:0]};

endmodule
